`timescale 1ns/1ps

module alu_test;

reg[31:0] i_datain, gr1, gr2;
wire[31:0] c, hi, lo;
wire zero, negative, overflow;

main test(i_datain, gr1, gr2, c, zero, negative, overflow, hi, lo);

initial
begin

$display("Instruction:op:func:ALUctr:ALUsrc:              gr1               :               gr2              :      imm       :shamt:                c               :   hi   :   lo   : zero : negative : overflow");
$monitor("   %h:%h: %h :  %h  :   %h  :%b:%b:%b:%b:%b:%h:%h:   %h  :     %h    :     %h",
i_datain, test.opcode, test.funct, test.aluctr, test.alusrc, gr1 , gr2, test.imm[15:0], test.shamt, c,
test.hi, test.lo, test.zero, test.negative, test.overflow);


//ADD: 1 + 8 = 9
#10 i_datain<=32'b000000_00011_00010_00001_00000_100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_1000;

//ADD: 2 + -2 = 0 zero
#10 i_datain<=32'b000000_00011_00010_00001_00000_100000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1110;

//ADD: -2 + -1 = -3 negative
#10 i_datain<=32'b000000_00011_00010_00001_00000_100000;
gr1<=32'b1111_1111_1111_1111_1111_1111_1111_1110;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

//ADD: -1 + -2147483648 = overflow
#10 i_datain<=32'b000000_00011_00010_00001_00000_100000;
gr1<=32'b1111_1111_1111_1111_1111_1111_1111_1111;
gr2<=32'b1000_0000_0000_0000_0000_0000_0000_0000;

//ADD: 2147483647 + 8 = overflow
#10 i_datain<=32'b000000_00011_00010_00001_00000_100000;
gr1<=32'b0111_1111_1111_1111_1111_1111_1111_1111;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_1000;



//ADDI: 7 + 8 = 15
#10 i_datain<=32'b001000_00011_00010_0000000000001000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0000;

//ADDI: 3 + -3 = 0 zero
#10 i_datain<=32'b001000_00011_00010_1111111111111101;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0000;

//ADDI: 1 + -64 = -63 negative
#10 i_datain<=32'b001000_00011_00010_1111111111000000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0000;

//ADDI: -2147483648 + -1 = overflow
#10 i_datain<=32'b001000_00011_00010_1111111111111111;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0000;



//ADDU: 2147483647 + 8 = 2147483655
#10 i_datain<=32'b000000_00011_00010_00001_00000_100001;
gr1<=32'b0111_1111_1111_1111_1111_1111_1111_1111;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_1000;



//ADDIU: 2147483647 + 8 = 2147483655
#10 i_datain<=32'b001001_00011_00010_0000000000001000;
gr1<=32'b0111_1111_1111_1111_1111_1111_1111_1111;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0000;



//SUB: 7 - 3 = 4
#10 i_datain<=32'b000000_00011_00010_00001_00000_100010;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

//SUB: 3 - 3 = 0 zero
#10 i_datain<=32'b000000_00011_00010_00001_00000_100010;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

//SUB: 3 - 7 = -4 negative
#10 i_datain<=32'b000000_00011_00010_00001_00000_100010;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0111;

//SUB: -2147483648 - 1 = overflow
#10 i_datain<=32'b000000_00011_00010_00001_00000_100010;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;



//SUBU: 2147483648 - 1 = 2147483647
#10 i_datain<=32'b000000_00011_00010_00001_00000_100011;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;



//MULT: 2 * 4 = 8
#10 i_datain<=32'b000000_00011_00010_00001_00000_011000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0100;

//MULT: 2 * 0 = 0 zero
#10 i_datain<=32'b000000_00011_00010_00001_00000_011000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0000;

//MULT: -2 * 4 = -8 negative
#10 i_datain<=32'b000000_00011_00010_00001_00000_011000;
gr1<=32'b1111_1111_1111_1111_1111_1111_1111_1110;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0100;

//MULT: 16777215 * 16777215 = 281474943156225
#10 i_datain<=32'b000000_00011_00010_00001_00000_011000;
gr1<=32'b0000_0000_1111_1111_1111_1111_1111_1111;
gr2<=32'b0000_0000_1111_1111_1111_1111_1111_1111;



//MULTU: 2147483649 * 1 = 2147483649
#10 i_datain<=32'b000000_00011_00010_00001_00000_011001;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;



//DIV: 8 / 3 = 2 ... 2
#10 i_datain<=32'b000000_00011_00010_00001_00000_011010;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_1000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

//DIV: 8 / -3 = -2 ... 2 negative
#10 i_datain<=32'b000000_00011_00010_00001_00000_011010;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_1000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1101;

//DIV: 2 / -3 = 0 ... 2 zero
#10 i_datain<=32'b000000_00011_00010_00001_00000_011010;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1101;

//DIV: -2147483648 / -1 = overflow
#10 i_datain<=32'b000000_00011_00010_00001_00000_011010;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;



//DIVU: 2147483648 / 1 = 2147483648 ... 0
#10 i_datain<=32'b000000_00011_00010_00001_00000_011011;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;



//AND: 1 & 2**32-1 = 1
#10 i_datain<=32'b000000_00011_00010_00001_00000_100100;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

//AND: 1 & 0 = 0
#10 i_datain<=32'b000000_00011_00010_00001_00000_100100;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0000;



//ANDI: 3 & 2**15+1 = 1
#10 i_datain<=32'b001100_00011_00010_1000000000000001;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0000;



//NOR: 4294967041 nor 241 = 14
#10 i_datain<=32'b000000_00011_00010_00001_00000_100111;
gr1<=32'b1111_1111_1111_1111_1111_1111_0000_0001;
gr2<=32'b0000_0000_0000_0000_0000_0000_1111_0001;

//NOR: 1 nor 2**32-1 = 0
#10 i_datain<=32'b000000_00011_00010_00001_00000_100111;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;



//OR: 11 | 4 = 15
#10 i_datain<=32'b000000_00011_00010_00001_00000_100101;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_1011;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0100;

//OR: 8 | 0 = 8
#10 i_datain<=32'b000000_00011_00010_00001_00000_100101;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_1000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0000;



//ORI: 3 & 2**15+5 = 2**15+7
#10 i_datain<=32'b001101_00011_00010_1000000000000101;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0000;




//XOR: 2**15 ^ 2**32-1 = 2*31-1
#10 i_datain<=32'b000000_00011_00010_00001_00000_100110;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;

//XOR: 3 ^ 7 = 4
#10 i_datain<=32'b000000_00011_00010_00001_00000_100110;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0111;



//XORI: 1 ^ 6 = 7
#10 i_datain<=32'b001110_00011_00010_0000000000000110;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0001;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;



//BEQ: 3 - 3 = 0 zero
#10 i_datain<=32'b000100_00011_00010_0000000000000111;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

//BEQ: 4 - 3 != 0
#10 i_datain<=32'b000100_00011_00010_0000000000000111;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;



//BNE: 3 - 3 = 0 zero
#10 i_datain<=32'b000101_00011_00010_0000000000000111;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;

//BNE: 4 - 3 != 0
#10 i_datain<=32'b000101_00011_00010_0000000000000111;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0100;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0011;



//SLT: 3 < 4 : 1
#10 i_datain<=32'b000000_00011_00010_00001_00000_101010;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0100;

//SLT: 7 < 4 : 0
#10 i_datain<=32'b000000_00011_00010_00001_00000_101010;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0100;

//SLT: 7 < -1 : 0
#10 i_datain<=32'b000000_00011_00010_00001_00000_101010;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;



//SLTI: 3 < 4 : 1
#10 i_datain<=32'b001010_00011_00010_0000000000000100;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0100;

//SLTI: 7 < -32768 : 0
#10 i_datain<=32'b001010_00011_00010_1000000000000000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0100;



//SLTIU: 7 < 2**15 : 1
#10 i_datain<=32'b001011_00011_00010_1000000000000000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;



//SLTU: 7 < 2**32-1 : 1
#10 i_datain<=32'b000000_00011_00010_00001_00000_101011;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0111;
gr2<=32'b1111_1111_1111_1111_1111_1111_1111_1111;



//LW: 8 + 4 = 12
#10 i_datain<=32'b100011_00011_00010_0000000000000100;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_1000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0100;



//SW: 2147483648 + -4 = 2147483644
#10 i_datain<=32'b100011_00011_00010_1111111111111100;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0100;



//SLL: 3 << 1 = 6 
#10 i_datain<=32'b000000_00011_00010_00001_00001_000000;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0111;

//SLL: 2**31 << 1 = 0
#10 i_datain<=32'b000000_00011_00010_00001_00001_000000;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0111;



//SLLV: 3 << 1 = 6 
#10 i_datain<=32'b000000_00011_00010_00001_00111_000100;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0011;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0001;



//SRL: 2**31 >> 21 = 2**10 = 1024
#10 i_datain<=32'b000000_00011_00010_00001_10101_000010;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0111;

//SRL: 2 >> 21 = 0
#10 i_datain<=32'b000000_00011_00010_00001_10101_000010;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_0010;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0111;



//SRLV: 9 >> 2 = 2
#10 i_datain<=32'b000000_00011_00010_00001_10101_000110;
gr1<=32'b0000_0000_0000_0000_0000_0000_0000_1001;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0010;



//SRA: -2147483648 >> 21 = -1024
#10 i_datain<=32'b000000_00011_00010_00001_10101_000011;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0000_0010;



//SRAV: -2147483648 >> 21 = -1024
#10 i_datain<=32'b000000_00011_00010_00001_00000_000111;
gr1<=32'b1000_0000_0000_0000_0000_0000_0000_0000;
gr2<=32'b0000_0000_0000_0000_0000_0000_0001_0101;



#10 $finish;
end
endmodule